module Not(s, r, q, qnot);

input a;
output y;

assign y = ~a;

endmodule
