// ----------------------------
// assign statements
//
// author: Tramy Nguyen
// ----------------------------

module simple_assign();
	
	reg a; 
	reg b;

	always begin 
		a = 1'b1;
		b = 1'b0;
	end
	
endmodule