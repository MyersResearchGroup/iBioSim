// ----------------------------
// An verilog module containing register declarations
//
// author: Tramy Nguyen
// ----------------------------

module registers();
	
	reg r1, r2, r3; 
	
endmodule