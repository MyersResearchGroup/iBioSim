// ----------------------------
// testing continuous assignments
//
// author: Tramy Nguyen
// ----------------------------

module contAssign(a, y);

  input a;
  output y;

assign y = ~a;

endmodule
