// ----------------------------
// if/else if/else statement
//
// author: Tramy Nguyen
// ----------------------------

module if_stmnt3();
	
	reg a, b; 

	always begin 
		if(a) begin
		end 
		else if(a) begin
		end
		else begin
		end
	end
	
endmodule