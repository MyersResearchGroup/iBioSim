// ----------------------------
// testing continuous assignments
//
// author: Tramy Nguyen
// ----------------------------

module contAssign4(a, b, y);

  input a;
  input b;
  output y;

assign y = a | b;
endmodule
